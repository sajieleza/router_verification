module router_top(clock,
                  resetn,
                  read_enb_0,
                  read_enb_1,
                  read_enb_2,
                  data_in,
                  pkt_valid,
                  busy,
                  error,
                  valid_out_0,
                  valid_out_1,
                  valid_out_2,
		  data_out_0,
                  data_out_1,
                  data_out_2);
input [7:0]data_in;
input clock,
      resetn,
      pkt_valid,
      read_enb_0,
      read_enb_1,
      read_enb_2;
output [7:0] data_out_0,data_out_1,data_out_2;
output busy,
       error,
       valid_out_0,
       valid_out_1,
       valid_out_2;

wire soft_reset_0,
     soft_reset_1,
     soft_reset_2,
     full_0,
     full_1,
     full_2,
     empty_0,
     empty_1,
     empty_2,
     fifo_full,
     detect_add,
     ld_state,
     laf_state,
     lfd_state,
     full_state,
     rst_int_reg,
     parity_done,
     low_pkt_valid,
     write_enb_reg;
wire [2:0]write_enb;
wire [7:0]data;

router_fifo FIFO_0(clock,resetn,write_enb[0],soft_reset_0,read_enb_0,data,lfd_state,empty_0,full_0,data_out_0);
router_fifo FIFO_1(clock,resetn,write_enb[1],soft_reset_1,read_enb_1,data,lfd_state,empty_1,full_1,data_out_1);
router_fifo FIFO_2(clock,resetn,write_enb[2],soft_reset_2,read_enb_2,data,lfd_state,empty_2,full_2,data_out_2);

router_reg REGISTER(clock,
                    resetn,
                    pkt_valid,
                    data_in,
                    fifo_full,
                    rst_int_reg,
                    detect_add,
                    ld_state,
                    laf_state,
                    full_state,
                    lfd_state,
                    parity_done,
                    low_pkt_valid,
                    error,
                    data);

router_sync SYNC(detect_add,
                   data_in[1:0],
                   write_enb_reg,
                   clock,
                   resetn,
                   valid_out_0,
                   valid_out_1,
                   valid_out_2,
                   read_enb_0,
                   read_enb_1,
                   read_enb_2,
                   write_enb,
                   fifo_full,
                   empty_0,
                   empty_1,
                   empty_2,
                   soft_reset_0,
                   soft_reset_1,
                   soft_reset_2,
                   full_0,
                   full_1,
                   full_2);

router_fsm FSM(clock,
                  resetn,
                  pkt_valid,
                  data_in[1:0],
                  fifo_full,
                  empty_0,
                  empty_1,
                  empty_2,
                  soft_reset_0,
                  soft_reset_1,
                  soft_reset_2,
		  parity_done,
                  low_pkt_valid,
                  write_enb_reg,
                  detect_add,
                  ld_state,
                  laf_state,
                  lfd_state,
                  full_state,
                  rst_int_reg,
                  busy);

endmodule
