//tb defns
